interface class DisplayElement;
    pure virtual local function void display();
endclass // DisplayElement
    
